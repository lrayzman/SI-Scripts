* 0;Circuit1.ckt

.CIRCUITNAME "Circuit1"
.rootnamemap 0;Circuit1
.namemap
W1=0;Circuit1;14
R1=0;Circuit1;2
L2=0;Circuit1;23
R3=0;Circuit1;4
L1=0;Circuit1;22
R2=0;Circuit1;3
C1=0;Circuit1;1
W2=0;Circuit1;21
C3=0;Circuit1;27
C4=0;Circuit1;28
C5=0;Circuit1;29
C2=0;Circuit1;24
.endnamemap
.stringparam syslib = "C:\Ansoft\DesignerSV2\DesignerSV2\syslib"
.stringparam userlib = "C:\Ansoft\DesignerSV2\DesignerSV2\userlib"
.stringparam personallib = "C:\Ansoft\DesignerSV2\MyProjects\PersonalLib"
.stringparam projectdir = "D:\Shared\Split_Deembedd"

*begin toplevel circuit

.SUB Microstrip MS(
+   H=6.6mil Er=3.50000000000000 TAND=0.0250000000000000 TANM=0 MSat=0 MRem=0
+MET1=1.72413800000000 T1=0.7mil)

MSTRL:14 net_65 net_6 W=10mil P=2500mil SUB=Microstrip
RES:2 0 net_6 R=150
IND:23 net_66 Port2 L=1nH 
RES:4 net_6 net_7 R=50
IND:22 Port1 net_65 L=1nH 
RES:3 0 net_7 R=150
CAP:1 net_6 net_7 C=10pF 
MSTRL:21 net_7 net_66 W=10mil P=2500mil SUB=Microstrip
CAP:27 0 net_65 C=0.5pF 
CAP:28 0 net_66 C=0.5pF 
CAP:29 0 Port2 C=0.5pF 
CAP:24 0 Port1 C=0.5pF 
PORT:Port2 Port2 0 PNUM=2 
PORT:Port1 Port1 0 PNUM=1 


*end toplevel circuit
.nwa:"NWA1"
+ F=LIN 0.01GHz 20GHz 0.01GHz
+ SWPORD = {F}
+ SolutionFile="C:\Ansoft\DesignerSV2\Temp\TestCase1.results\Circuit1_NWA1_105_U1_Circuit1_107_0\Circuit1_NWA1_105_U1_Circuit1_107_0.sol"

.end
