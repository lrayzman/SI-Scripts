* 176;E2E.ckt

.CIRCUITNAME "E2E"
.rootnamemap 176;E2E
.namemap
C1=176;E2E;1
R1=176;E2E;2
R2=176;E2E;3
R3=176;E2E;4
W1=176;E2E;14
W2=176;E2E;21
L1=176;E2E;22
L2=176;E2E;23
C2=176;E2E;24
C3=176;E2E;27
C4=176;E2E;28
C5=176;E2E;29
.endnamemap
.stringparam syslib = "C:\Ansoft\DesignerSV2\DesignerSV2\syslib"
.stringparam userlib = "C:\Ansoft\DesignerSV2\DesignerSV2\userlib"
.stringparam personallib = "C:\Ansoft\DesignerSV2\MyProjects\PersonalLib"
.stringparam projectdir = "D:\Shared\Split_Deembedd"

*begin toplevel circuit

.SUB Microstrip MS(
+   H=6.6mil Er=3.50000000000000 TAND=0.0250000000000000 TANM=0 MSat=0 MRem=0
+MET1=1.72413800000000 T1=0.7mil)

CAP:1 net_6 net_7 C=15pF 
RES:2 0 net_6 R=1000
RES:3 0 net_7 R=1000
RES:4 net_6 net_7 R=50
MSTRL:14 net_65 net_6 W=10mil P=2500mil SUB=Microstrip
MSTRL:21 net_7 net_66 W=10mil P=2500mil SUB=Microstrip
IND:22 Port1 net_65 L=0.25nH 
IND:23 net_66 Port2 L=0.25nH 
CAP:24 0 Port1 C=0.25pF 
CAP:27 0 net_65 C=0.25pF 
CAP:28 0 net_66 C=0.25pF 
CAP:29 0 Port2 C=0.25pF 
PORT:Port1 Port1 0 PNUM=1 
PORT:Port2 Port2 0 PNUM=2 rz=50Ohm iz=0Ohm 


*end toplevel circuit
.nwa:"NWA1"
+ F=LIN 0.01GHz 20GHz 0.01GHz
+ SWPORD = {F}
+ SolutionFile="C:\Ansoft\DesignerSV2\Temp\TestCase1.results\E2E_NWA1_105_U4_E2E_0_73\E2E_NWA1_105_U4_E2E_0_73.sol"

.end
